(a+(b))*(c)/(d)+((func(func2(a+(b*c+func3(1))))+c)*d);